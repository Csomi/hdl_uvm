
package my_pkg;
	`include "uvm_macros.svh"
	import uvm_pkg::*;
	`include "my_env.svh"
	`include "my_first_test.svh"
endpackage: my_pkg
